module exe_initiator  ( output logic base_addr,
						output logic pdp_mem_opcode,
						output logic pdp_op7_opcode,
						input stall,
						input PC_value);
						
						
